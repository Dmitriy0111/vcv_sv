/*
*  File            :   keyboard_pkg.sv
*  Autor           :   Vlasov D.V
*  Data            :   15.05.2020
*  Language        :   SystemVerilog
*  Description     :   This is keyboard package
*  Copyright(c)    :   2019-2020 Vlasov D.V
*/

package keyboard_pkg;

    `include    "keyboard_c.sv"

endpackage: keyboard_pkg
